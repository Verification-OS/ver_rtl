
// NOTE: User is free to add more cover properties in this file that is included FV_cov.sv.
