
`protect

`ifndef _FV_SI_LATENCIES_DUT_SVH
`define _FV_SI_LATENCIES_DUT_SVH

`define FV_SI_LATENCY_ALU  (6 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_ADD  `FV_SI_LATENCY_ALU
`define FV_SI_LATENCY_SUB  `FV_SI_LATENCY_ALU
`define FV_SI_LATENCY_SLL  `FV_SI_LATENCY_ALU
`define FV_SI_LATENCY_SLT  `FV_SI_LATENCY_ALU
`define FV_SI_LATENCY_SLTU `FV_SI_LATENCY_ALU
`define FV_SI_LATENCY_XOR  `FV_SI_LATENCY_ALU
`define FV_SI_LATENCY_SRL  `FV_SI_LATENCY_ALU
`define FV_SI_LATENCY_SRA  `FV_SI_LATENCY_ALU
`define FV_SI_LATENCY_OR   `FV_SI_LATENCY_ALU
`define FV_SI_LATENCY_AND  `FV_SI_LATENCY_ALU

`define FV_SI_LATENCY_LUI   `FV_SI_LATENCY_ALU
`define FV_SI_LATENCY_AUIPC `FV_SI_LATENCY_ALU

`define FV_SI_LATENCY_MUL_ALL (8 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_MUL    `FV_SI_LATENCY_MUL_ALL
`define FV_SI_LATENCY_MULH   `FV_SI_LATENCY_MUL_ALL
`define FV_SI_LATENCY_MULHSU `FV_SI_LATENCY_MUL_ALL
`define FV_SI_LATENCY_MULHU  `FV_SI_LATENCY_MUL_ALL

`define FV_SI_LATENCY_DIV_ALL (38+ `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_DIV  `FV_SI_LATENCY_DIV_ALL
`define FV_SI_LATENCY_DIVU `FV_SI_LATENCY_DIV_ALL
`define FV_SI_LATENCY_REM  `FV_SI_LATENCY_DIV_ALL
`define FV_SI_LATENCY_REMU `FV_SI_LATENCY_DIV_ALL

`define FV_SI_LATENCY_LB (14 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_LH (14 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_LW (14 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_LD (14 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_LBU (14 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_LHU (14 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_LWU (14 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_SB (11 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_SH (11 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_SW (11 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_SD (11 + `FV_SI_FE_PIPE_DELAY)

`define FV_SI_LATENCY_JMP (6 + `FV_SI_FE_PIPE_DELAY)

`define FV_SI_LATENCY_AMOW (18 + `FV_SI_FE_PIPE_DELAY)
`define FV_SI_LATENCY_AMOD (18 + `FV_SI_FE_PIPE_DELAY)

`endif //  `ifndef _FV_SI_LATENCIES_DUT_SVH

`endprotect
